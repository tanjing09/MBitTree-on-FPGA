`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2021/09/02 11:41:06
// Design Name: 
// Module Name: testbench_sa
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module testbench_sa 
(
    );
    
    
    reg clk;
    reg RSTn;
    reg [104-1:0] packet_in1;
    reg           data_valid_in1;
    reg [104-1:0] packet_in2;
    reg           data_valid_in2;
    
    wire [14-1:0] rule_id1;
    wire [14-1:0] rule_id2;
    wire          data_valid_out1;
    wire          data_valid_out2;
    wire          action_valid1;
    wire          action_valid2;
    
    initial begin
        clk = 1'b1;
        forever begin
            #2 clk = ~clk;
        end
    end
    
    initial begin
        RSTn = 1'b0;
        #20 RSTn = 1'b1;
    end
    
    initial begin
        packet_in1 = 104'bX;
        packet_in2 = 104'bX;
        data_valid_in1 = 1'b0;
        data_valid_in2 = 1'b0;
        #40
        //3817,4562
        packet_in1 = 104'b00000001_0000000000000000_0000000000000000_01000000000000000000000000000000_00010110000101010000001011000001;
        packet_in2 = 104'b00000001_1111111111111111_1111111111111111_10000000000000000000000000000000_00000110101000100001000000000000;
        data_valid_in1 = 1'b1;
        data_valid_in2 = 1'b1;
        #4
        //4457,4635
        packet_in1 = 104'b00000001_1111111111111111_1111111111111111_10000000000000000000000000000000_00100010100101000001100011100000;
        packet_in2 = 104'b00000001_1111111111111111_1111111111111111_11111111111111111111111111111111_00111010001011000101101110101011;
        data_valid_in1 = 1'b1;
        data_valid_in2 = 1'b1;
        #4
        //4480,4444
        packet_in1 = 104'b00000001_0000000000000000_0000000000000000_11111111111111111111111111111111_00010111010110010000001001100000;
        packet_in2 = 104'b00000001_0000000000000000_0000000000000000_11111111111111111111111111111111_00111001010001111000101111100010;
        data_valid_in1 = 1'b1;
        data_valid_in2 = 1'b1;
        #4
        //6764, 6826
        packet_in1 = 104'b00000001_0000000000000000_1111111111111111_00000000000000000000000000000000_00100110111111101101011100000011;
        packet_in2 = 104'b00000001_1111111111111111_1111111111111111_00000000000000000000000000000000_00001100110011011000110001000010;
        data_valid_in1 = 1'b1;
        data_valid_in2 = 1'b1;
        #4
        //4634, 7385
        packet_in1 = 104'b00000001_0000000000000000_0000000000000000_11111111111111111111111111111111_00111010000011001100011001000011;
        packet_in2 = 104'b00000000_0000000000000000_1111111111111111_01000000000000000000000000000000_00110100111011010100011100101011;
        data_valid_in1 = 1'b1;
        data_valid_in2 = 1'b1;
        #4
        //3806, 4667
        packet_in1 = 104'b00000001_1111111111111111_0000000000000000_01000000000000000000000000000000_00110011011010000000011111101001;
        packet_in2 = 104'b00000001_0000000000000000_0000000000000000_00000000000000000000000000000000_00101111010101000101111000101010;
        data_valid_in1 = 1'b1;
        data_valid_in2 = 1'b1;
        #4
        //4474, 4449
        packet_in1 = 104'b00000001_0000000000000000_1111111111111111_10000000000000000000000000000000_00010001111010111001111100001010;
        packet_in2 = 104'b00000001_1111111111111111_1111111111111111_10000000000000000000000000000000_00110101101010011001110101000000;
        data_valid_in1 = 1'b1;
        data_valid_in2 = 1'b1;
        #4
        //4696,3809
        packet_in1 = 104'b00000001111111111111111111111111111111110000000000000000000000000000000000000010100011010000100100010000;
        packet_in2 = 104'b00000001111111111111111111111111111111110100000000000000000000000000000000101010011010111100101001111000;
        data_valid_in1 = 1'b1;
        data_valid_in2 = 1'b1;
        #4
        //6795, 4529
        packet_in1 = 104'b00000001111111111111111111111111111111110000000000000000000000000000000000011100110000000001001001011010;
        packet_in2 = 104'b00000001111111111111111100000000000000001111111111111111111111111111111100111100101110111101101101011000;
        data_valid_in1 = 1'b1;
        data_valid_in2 = 1'b1;
        #4
        //4491, 3802
        packet_in1 = 104'b00000001111111111111111111111111111111111000000000000000000000000000000000000101010000011000000111011011;
        packet_in2 = 104'b00000001000000000000000011111111111111110111111111111111111111111111111100111101001101111101000011011011;
        data_valid_in1 = 1'b1;
        data_valid_in2 = 1'b1;
        #4
        packet_in1 = 104'b0;
        packet_in2 = 104'b0;
        data_valid_in1 = 1'b0;
        data_valid_in2 = 1'b0;
    end
    
    pipeline_SA pipeline_SA_inst(
        .clk(clk),
        .RSTn(RSTn),
    
        //dual port
        .packet_in1 (packet_in1),
        .packet_in2 (packet_in2),
        .data_valid_in1 (data_valid_in1),
        .data_valid_in2 (data_valid_in2),
        
        .rule_id1 (rule_id1),
        .rule_id2 (rule_id2),
        .data_valid_out1 (data_valid_out1),
        .data_valid_out2 (data_valid_out2),
        .action_valid1 (action_valid1),
        .action_valid2 (action_valid2)    
    );
    
endmodule
